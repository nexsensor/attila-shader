//Author  :Alex Zhang (cgalexzhang@sina.com)
//Date    :01-05-2020
//Comment : a subset of Attila Shader Instructions
module attila_shader (
input  gclk,
input  resetn,

);



endmoudle 
